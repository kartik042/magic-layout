magic
tech scmos
timestamp 1461907805
<< nwell >>
rect -40 8 70 30
rect 115 8 225 30
rect -7 -69 33 -53
rect 137 -57 177 -41
rect 201 -70 241 -54
<< polysilicon >>
rect 2 20 54 22
rect -28 14 -26 16
rect -6 14 -4 16
rect 2 14 4 20
rect 24 14 26 16
rect 32 14 34 16
rect 52 14 54 20
rect 157 20 209 22
rect 127 14 129 16
rect 149 14 151 16
rect 157 14 159 20
rect 179 14 181 16
rect 187 14 189 16
rect 207 14 209 20
rect -28 -18 -26 10
rect -6 2 -4 10
rect -16 0 -4 2
rect -28 -24 -26 -22
rect -16 -26 -14 0
rect 2 -2 4 10
rect -8 -4 4 -2
rect -8 -14 -6 -4
rect 24 -10 26 10
rect 6 -12 26 -10
rect -8 -16 -4 -14
rect -6 -18 -4 -16
rect 6 -18 8 -12
rect 24 -18 26 -16
rect 32 -18 34 10
rect 52 -18 54 10
rect 127 -18 129 10
rect 149 2 151 10
rect 139 0 151 2
rect -6 -24 -4 -22
rect 6 -24 8 -22
rect 24 -26 26 -22
rect 32 -24 34 -22
rect 52 -24 54 -22
rect 127 -24 129 -22
rect -16 -28 26 -26
rect 139 -26 141 0
rect 157 -2 159 10
rect 147 -4 159 -2
rect 147 -14 149 -4
rect 179 -10 181 10
rect 161 -12 181 -10
rect 147 -16 151 -14
rect 149 -18 151 -16
rect 161 -18 163 -12
rect 179 -18 181 -16
rect 187 -18 189 10
rect 207 -18 209 10
rect 149 -24 151 -22
rect 161 -24 163 -22
rect 179 -26 181 -22
rect 187 -24 189 -22
rect 207 -24 209 -22
rect 139 -28 181 -26
rect 151 -51 153 -49
rect 161 -51 163 -49
rect 7 -63 9 -61
rect 17 -63 19 -61
rect 7 -93 9 -67
rect 17 -93 19 -67
rect 151 -81 153 -55
rect 161 -81 163 -55
rect 215 -64 217 -62
rect 225 -64 227 -62
rect 151 -87 153 -85
rect 161 -87 163 -85
rect 215 -94 217 -68
rect 225 -94 227 -68
rect 7 -99 9 -97
rect 17 -99 19 -97
rect 215 -100 217 -98
rect 225 -100 227 -98
<< ndiffusion >>
rect -32 -22 -28 -18
rect -26 -22 -22 -18
rect -8 -22 -6 -18
rect -4 -22 6 -18
rect 8 -22 10 -18
rect 22 -22 24 -18
rect 26 -22 32 -18
rect 34 -22 36 -18
rect 48 -22 52 -18
rect 54 -22 58 -18
rect 123 -22 127 -18
rect 129 -22 133 -18
rect 147 -22 149 -18
rect 151 -22 161 -18
rect 163 -22 165 -18
rect 177 -22 179 -18
rect 181 -22 187 -18
rect 189 -22 191 -18
rect 203 -22 207 -18
rect 209 -22 213 -18
rect 141 -85 143 -81
rect 147 -85 151 -81
rect 153 -85 161 -81
rect 163 -85 167 -81
rect 171 -85 173 -81
rect -3 -97 -1 -93
rect 3 -97 7 -93
rect 9 -97 17 -93
rect 19 -97 23 -93
rect 27 -97 29 -93
rect 205 -98 207 -94
rect 211 -98 215 -94
rect 217 -98 225 -94
rect 227 -98 231 -94
rect 235 -98 237 -94
<< pdiffusion >>
rect -32 10 -28 14
rect -26 10 -22 14
rect -8 10 -6 14
rect -4 10 2 14
rect 4 10 10 14
rect 22 10 24 14
rect 26 10 32 14
rect 34 10 36 14
rect 48 10 52 14
rect 54 10 58 14
rect 123 10 127 14
rect 129 10 133 14
rect 147 10 149 14
rect 151 10 157 14
rect 159 10 165 14
rect 177 10 179 14
rect 181 10 187 14
rect 189 10 191 14
rect 203 10 207 14
rect 209 10 213 14
rect 141 -55 143 -51
rect 147 -55 151 -51
rect 153 -55 155 -51
rect 159 -55 161 -51
rect 163 -55 167 -51
rect 171 -55 173 -51
rect -3 -67 -1 -63
rect 3 -67 7 -63
rect 9 -67 11 -63
rect 15 -67 17 -63
rect 19 -67 23 -63
rect 27 -67 29 -63
rect 205 -68 207 -64
rect 211 -68 215 -64
rect 217 -68 219 -64
rect 223 -68 225 -64
rect 227 -68 231 -64
rect 235 -68 237 -64
<< metal1 >>
rect -36 24 -20 28
rect -16 24 14 28
rect 18 24 48 28
rect 52 24 66 28
rect 119 24 135 28
rect 139 24 169 28
rect 173 24 203 28
rect 207 24 221 28
rect -36 14 -32 24
rect -12 14 -8 24
rect 36 14 40 24
rect 58 14 62 24
rect -22 6 -18 10
rect -22 2 -10 6
rect -48 -6 -32 -2
rect -48 -73 -44 -6
rect -40 -10 -36 -6
rect -22 -18 -18 2
rect 0 -10 6 -8
rect 0 -12 2 -10
rect 10 -18 14 10
rect 119 14 123 24
rect 143 14 147 24
rect 191 14 195 24
rect 213 14 217 24
rect 18 -18 22 10
rect 44 -8 48 10
rect 133 6 137 10
rect 62 2 110 6
rect 38 -12 48 -8
rect 106 -2 110 2
rect 133 2 145 6
rect 106 -6 123 -2
rect 44 -18 48 -12
rect 58 -14 74 -10
rect -36 -28 -32 -22
rect -12 -28 -8 -22
rect 36 -28 40 -22
rect 58 -28 62 -22
rect -36 -32 -22 -28
rect -18 -32 28 -28
rect 32 -32 46 -28
rect 50 -32 66 -28
rect -5 -59 -1 -55
rect 3 -59 11 -55
rect 15 -59 23 -55
rect 27 -59 31 -55
rect -1 -63 3 -59
rect 23 -63 27 -59
rect 11 -73 15 -67
rect -48 -77 3 -73
rect 11 -77 27 -73
rect -12 -87 13 -83
rect 23 -84 27 -77
rect -12 -108 -8 -87
rect 23 -93 27 -88
rect -1 -101 3 -97
rect -5 -105 -1 -101
rect 3 -105 12 -101
rect 16 -105 23 -101
rect 27 -105 31 -101
rect 70 -108 74 -14
rect 106 -71 110 -6
rect 115 -10 119 -6
rect 133 -18 137 2
rect 155 -10 161 -8
rect 155 -12 157 -10
rect 165 -18 169 10
rect 173 -18 177 10
rect 199 -8 203 10
rect 218 2 224 6
rect 193 -12 203 -8
rect 199 -18 203 -12
rect 213 -14 230 -10
rect 119 -28 123 -22
rect 143 -28 147 -22
rect 191 -28 195 -22
rect 213 -28 217 -22
rect 119 -32 133 -28
rect 137 -32 183 -28
rect 187 -32 201 -28
rect 205 -32 221 -28
rect 226 -36 230 -14
rect 128 -40 230 -36
rect 128 -61 132 -40
rect 139 -47 143 -43
rect 147 -47 155 -43
rect 159 -47 167 -43
rect 171 -47 175 -43
rect 143 -51 147 -47
rect 167 -51 171 -47
rect 155 -61 159 -55
rect 203 -60 207 -56
rect 211 -60 219 -56
rect 223 -60 231 -56
rect 235 -60 239 -56
rect 128 -65 147 -61
rect 155 -65 171 -61
rect 106 -75 157 -71
rect 167 -74 171 -65
rect 207 -64 211 -60
rect 231 -64 235 -60
rect 219 -74 223 -68
rect 167 -78 211 -74
rect 219 -78 235 -74
rect 167 -81 171 -78
rect 143 -89 147 -85
rect 204 -88 221 -84
rect 139 -93 143 -89
rect 147 -93 155 -89
rect 159 -93 167 -89
rect 171 -93 175 -89
rect 231 -94 235 -78
rect 207 -102 211 -98
rect 203 -106 207 -102
rect 211 -106 219 -102
rect 223 -106 231 -102
rect 235 -106 239 -102
rect -12 -112 74 -108
<< metal2 >>
rect 18 2 58 6
rect 173 2 214 6
rect -12 -10 -4 -8
rect -36 -12 -4 -10
rect 143 -10 151 -8
rect -36 -14 -8 -12
rect 119 -12 151 -10
rect 119 -14 147 -12
rect 27 -88 110 -84
rect 106 -98 110 -88
rect 192 -88 200 -84
rect 192 -98 196 -88
rect 106 -102 196 -98
<< ntransistor >>
rect -28 -22 -26 -18
rect -6 -22 -4 -18
rect 6 -22 8 -18
rect 24 -22 26 -18
rect 32 -22 34 -18
rect 52 -22 54 -18
rect 127 -22 129 -18
rect 149 -22 151 -18
rect 161 -22 163 -18
rect 179 -22 181 -18
rect 187 -22 189 -18
rect 207 -22 209 -18
rect 151 -85 153 -81
rect 161 -85 163 -81
rect 7 -97 9 -93
rect 17 -97 19 -93
rect 215 -98 217 -94
rect 225 -98 227 -94
<< ptransistor >>
rect -28 10 -26 14
rect -6 10 -4 14
rect 2 10 4 14
rect 24 10 26 14
rect 32 10 34 14
rect 52 10 54 14
rect 127 10 129 14
rect 149 10 151 14
rect 157 10 159 14
rect 179 10 181 14
rect 187 10 189 14
rect 207 10 209 14
rect 151 -55 153 -51
rect 161 -55 163 -51
rect 7 -67 9 -63
rect 17 -67 19 -63
rect 215 -68 217 -64
rect 225 -68 227 -64
<< polycontact >>
rect -32 -6 -28 -2
rect -10 2 -6 6
rect 2 -14 6 -10
rect 34 -12 38 -8
rect 123 -6 127 -2
rect 54 -14 58 -10
rect 145 2 149 6
rect 157 -14 161 -10
rect 189 -12 193 -8
rect 209 -14 213 -10
rect 147 -65 151 -61
rect 3 -77 7 -73
rect 13 -87 17 -83
rect 157 -75 161 -71
rect 211 -78 215 -74
rect 221 -88 225 -84
<< ndcontact >>
rect -36 -22 -32 -18
rect -22 -22 -18 -18
rect -12 -22 -8 -18
rect 10 -22 14 -18
rect 18 -22 22 -18
rect 36 -22 40 -18
rect 44 -22 48 -18
rect 58 -22 62 -18
rect 119 -22 123 -18
rect 133 -22 137 -18
rect 143 -22 147 -18
rect 165 -22 169 -18
rect 173 -22 177 -18
rect 191 -22 195 -18
rect 199 -22 203 -18
rect 213 -22 217 -18
rect 143 -85 147 -81
rect 167 -85 171 -81
rect -1 -97 3 -93
rect 23 -97 27 -93
rect 207 -98 211 -94
rect 231 -98 235 -94
<< pdcontact >>
rect -36 10 -32 14
rect -22 10 -18 14
rect -12 10 -8 14
rect 10 10 14 14
rect 18 10 22 14
rect 36 10 40 14
rect 44 10 48 14
rect 58 10 62 14
rect 119 10 123 14
rect 133 10 137 14
rect 143 10 147 14
rect 165 10 169 14
rect 173 10 177 14
rect 191 10 195 14
rect 199 10 203 14
rect 213 10 217 14
rect 143 -55 147 -51
rect 155 -55 159 -51
rect 167 -55 171 -51
rect -1 -67 3 -63
rect 11 -67 15 -63
rect 23 -67 27 -63
rect 207 -68 211 -64
rect 219 -68 223 -64
rect 231 -68 235 -64
<< m2contact >>
rect -40 -14 -36 -10
rect -4 -12 0 -8
rect 14 2 18 6
rect 58 2 62 6
rect 23 -88 27 -84
rect 115 -14 119 -10
rect 151 -12 155 -8
rect 169 2 173 6
rect 214 2 218 6
rect 200 -88 204 -84
<< psubstratepcontact >>
rect -22 -32 -18 -28
rect 28 -32 32 -28
rect 46 -32 50 -28
rect 133 -32 137 -28
rect 183 -32 187 -28
rect 201 -32 205 -28
rect 143 -93 147 -89
rect 155 -93 159 -89
rect 167 -93 171 -89
rect -1 -105 3 -101
rect 12 -105 16 -101
rect 23 -105 27 -101
rect 207 -106 211 -102
rect 219 -106 223 -102
rect 231 -106 235 -102
<< nsubstratencontact >>
rect -20 24 -16 28
rect 14 24 18 28
rect 48 24 52 28
rect 135 24 139 28
rect 169 24 173 28
rect 203 24 207 28
rect 143 -47 147 -43
rect 155 -47 159 -43
rect 167 -47 171 -43
rect -1 -59 3 -55
rect 11 -59 15 -55
rect 23 -59 27 -55
rect 207 -60 211 -56
rect 219 -60 223 -56
rect 231 -60 235 -56
<< labels >>
rlabel polycontact -30 -5 -28 -3 1 A
rlabel polycontact 54 -13 56 -11 1 B
rlabel metal1 4 25 6 27 5 VDD
rlabel metal1 8 -31 10 -29 1 GND
rlabel metal1 159 25 161 27 5 VDD
rlabel metal1 163 -31 165 -29 1 GND
rlabel nsubstratencontact 156 -46 158 -44 1 VDD
rlabel psubstratepcontact 156 -92 158 -90 1 GND
rlabel nsubstratencontact 12 -58 14 -56 1 VDD
rlabel psubstratepcontact 12 -104 14 -102 1 GND
rlabel nsubstratencontact 220 -59 222 -57 1 VDD
rlabel psubstratepcontact 220 -105 222 -103 1 GND
rlabel metal1 129 -39 131 -37 1 Cin
rlabel metal1 221 3 223 5 1 Sum
rlabel metal1 232 -77 234 -75 1 Cout
<< end >>
