magic
tech scmos
timestamp 1459893001
<< polysilicon >>
rect -8 44 -4 48
rect 14 44 18 48
rect -8 -26 -4 32
rect 14 -26 18 32
rect -8 -40 -4 -36
rect 14 -40 18 -36
<< ndiffusion >>
rect -22 -30 -8 -26
rect -22 -36 -20 -30
rect -14 -36 -8 -30
rect -4 -36 14 -26
rect 18 -32 28 -26
rect 18 -36 34 -32
<< pdiffusion >>
rect -22 38 -18 44
rect -12 38 -8 44
rect -22 32 -8 38
rect -4 38 14 44
rect -4 32 2 38
rect 8 32 14 38
rect 18 38 22 44
rect 28 38 32 44
rect 18 32 32 38
<< metal1 >>
rect -22 58 32 68
rect -18 44 -12 58
rect 22 44 28 58
rect 2 20 8 32
rect -20 14 -12 18
rect 2 14 44 20
rect -20 -8 18 -4
rect 28 -26 34 14
rect -20 -48 -14 -36
rect -22 -56 34 -48
<< ntransistor >>
rect -8 -36 -4 -26
rect 14 -36 18 -26
<< ptransistor >>
rect -8 32 -4 44
rect 14 32 18 44
<< polycontact >>
rect -12 14 -8 18
rect 18 -8 22 -4
<< ndcontact >>
rect -20 -36 -14 -30
rect 28 -32 34 -26
<< pdcontact >>
rect -18 38 -12 44
rect 2 32 8 38
rect 22 38 28 44
<< labels >>
rlabel metal1 -20 14 -8 18 1 A
rlabel metal1 -20 -8 -8 -4 1 B
rlabel metal1 -22 -56 34 -48 1 GND
rlabel metal1 -22 58 32 68 5 VDD
rlabel metal1 34 14 44 20 7 Y
<< end >>
