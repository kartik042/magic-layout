magic
tech scmos
timestamp 1461965142
<< nwell >>
rect -40 8 70 30
rect 115 8 225 30
rect 264 9 374 31
rect 419 9 529 31
rect 568 9 678 31
rect 723 9 833 31
rect 873 9 983 31
rect 1028 9 1138 31
rect -7 -69 33 -53
rect 137 -57 177 -41
rect 201 -70 241 -54
rect 297 -68 337 -52
rect 441 -56 481 -40
rect 505 -69 545 -53
rect 601 -68 641 -52
rect 745 -56 785 -40
rect 809 -69 849 -53
rect 906 -68 946 -52
rect 1050 -56 1090 -40
rect 1114 -69 1154 -53
<< polysilicon >>
rect 2 20 54 22
rect -28 14 -26 16
rect -6 14 -4 16
rect 2 14 4 20
rect 24 14 26 16
rect 32 14 34 16
rect 52 14 54 20
rect 157 20 209 22
rect 127 14 129 16
rect 149 14 151 16
rect 157 14 159 20
rect 179 14 181 16
rect 187 14 189 16
rect 207 14 209 20
rect 306 21 358 23
rect 276 15 278 17
rect 298 15 300 17
rect 306 15 308 21
rect 328 15 330 17
rect 336 15 338 17
rect 356 15 358 21
rect 461 21 513 23
rect 431 15 433 17
rect 453 15 455 17
rect 461 15 463 21
rect 483 15 485 17
rect 491 15 493 17
rect 511 15 513 21
rect 610 21 662 23
rect 580 15 582 17
rect 602 15 604 17
rect 610 15 612 21
rect 632 15 634 17
rect 640 15 642 17
rect 660 15 662 21
rect 765 21 817 23
rect 735 15 737 17
rect 757 15 759 17
rect 765 15 767 21
rect 787 15 789 17
rect 795 15 797 17
rect 815 15 817 21
rect 915 21 967 23
rect 885 15 887 17
rect 907 15 909 17
rect 915 15 917 21
rect 937 15 939 17
rect 945 15 947 17
rect 965 15 967 21
rect 1070 21 1122 23
rect 1040 15 1042 17
rect 1062 15 1064 17
rect 1070 15 1072 21
rect 1092 15 1094 17
rect 1100 15 1102 17
rect 1120 15 1122 21
rect -28 -18 -26 10
rect -6 2 -4 10
rect -16 0 -4 2
rect -28 -24 -26 -22
rect -16 -26 -14 0
rect 2 -2 4 10
rect -8 -4 4 -2
rect -8 -14 -6 -4
rect 24 -10 26 10
rect 6 -12 26 -10
rect -8 -16 -4 -14
rect -6 -18 -4 -16
rect 6 -18 8 -12
rect 24 -18 26 -16
rect 32 -18 34 10
rect 52 -18 54 10
rect 127 -18 129 10
rect 149 2 151 10
rect 139 0 151 2
rect -6 -24 -4 -22
rect 6 -24 8 -22
rect 24 -26 26 -22
rect 32 -24 34 -22
rect 52 -24 54 -22
rect 127 -24 129 -22
rect -16 -28 26 -26
rect 139 -26 141 0
rect 157 -2 159 10
rect 147 -4 159 -2
rect 147 -14 149 -4
rect 179 -10 181 10
rect 161 -12 181 -10
rect 147 -16 151 -14
rect 149 -18 151 -16
rect 161 -18 163 -12
rect 179 -18 181 -16
rect 187 -18 189 10
rect 207 -18 209 10
rect 276 -17 278 11
rect 298 3 300 11
rect 288 1 300 3
rect 149 -24 151 -22
rect 161 -24 163 -22
rect 179 -26 181 -22
rect 187 -24 189 -22
rect 207 -24 209 -22
rect 276 -23 278 -21
rect 139 -28 181 -26
rect 288 -25 290 1
rect 306 -1 308 11
rect 296 -3 308 -1
rect 296 -13 298 -3
rect 328 -9 330 11
rect 310 -11 330 -9
rect 296 -15 300 -13
rect 298 -17 300 -15
rect 310 -17 312 -11
rect 328 -17 330 -15
rect 336 -17 338 11
rect 356 -17 358 11
rect 431 -17 433 11
rect 453 3 455 11
rect 443 1 455 3
rect 298 -23 300 -21
rect 310 -23 312 -21
rect 328 -25 330 -21
rect 336 -23 338 -21
rect 356 -23 358 -21
rect 431 -23 433 -21
rect 288 -27 330 -25
rect 443 -25 445 1
rect 461 -1 463 11
rect 451 -3 463 -1
rect 451 -13 453 -3
rect 483 -9 485 11
rect 465 -11 485 -9
rect 451 -15 455 -13
rect 453 -17 455 -15
rect 465 -17 467 -11
rect 483 -17 485 -15
rect 491 -17 493 11
rect 511 -17 513 11
rect 580 -17 582 11
rect 602 3 604 11
rect 592 1 604 3
rect 453 -23 455 -21
rect 465 -23 467 -21
rect 483 -25 485 -21
rect 491 -23 493 -21
rect 511 -23 513 -21
rect 580 -23 582 -21
rect 443 -27 485 -25
rect 592 -25 594 1
rect 610 -1 612 11
rect 600 -3 612 -1
rect 600 -13 602 -3
rect 632 -9 634 11
rect 614 -11 634 -9
rect 600 -15 604 -13
rect 602 -17 604 -15
rect 614 -17 616 -11
rect 632 -17 634 -15
rect 640 -17 642 11
rect 660 -17 662 11
rect 735 -17 737 11
rect 757 3 759 11
rect 747 1 759 3
rect 602 -23 604 -21
rect 614 -23 616 -21
rect 632 -25 634 -21
rect 640 -23 642 -21
rect 660 -23 662 -21
rect 735 -23 737 -21
rect 592 -27 634 -25
rect 747 -25 749 1
rect 765 -1 767 11
rect 755 -3 767 -1
rect 755 -13 757 -3
rect 787 -9 789 11
rect 769 -11 789 -9
rect 755 -15 759 -13
rect 757 -17 759 -15
rect 769 -17 771 -11
rect 787 -17 789 -15
rect 795 -17 797 11
rect 815 -17 817 11
rect 885 -17 887 11
rect 907 3 909 11
rect 897 1 909 3
rect 757 -23 759 -21
rect 769 -23 771 -21
rect 787 -25 789 -21
rect 795 -23 797 -21
rect 815 -23 817 -21
rect 885 -23 887 -21
rect 747 -27 789 -25
rect 897 -25 899 1
rect 915 -1 917 11
rect 905 -3 917 -1
rect 905 -13 907 -3
rect 937 -9 939 11
rect 919 -11 939 -9
rect 905 -15 909 -13
rect 907 -17 909 -15
rect 919 -17 921 -11
rect 937 -17 939 -15
rect 945 -17 947 11
rect 965 -17 967 11
rect 1040 -17 1042 11
rect 1062 3 1064 11
rect 1052 1 1064 3
rect 907 -23 909 -21
rect 919 -23 921 -21
rect 937 -25 939 -21
rect 945 -23 947 -21
rect 965 -23 967 -21
rect 1040 -23 1042 -21
rect 897 -27 939 -25
rect 1052 -25 1054 1
rect 1070 -1 1072 11
rect 1060 -3 1072 -1
rect 1060 -13 1062 -3
rect 1092 -9 1094 11
rect 1074 -11 1094 -9
rect 1060 -15 1064 -13
rect 1062 -17 1064 -15
rect 1074 -17 1076 -11
rect 1092 -17 1094 -15
rect 1100 -17 1102 11
rect 1120 -17 1122 11
rect 1062 -23 1064 -21
rect 1074 -23 1076 -21
rect 1092 -25 1094 -21
rect 1100 -23 1102 -21
rect 1120 -23 1122 -21
rect 1052 -27 1094 -25
rect 151 -51 153 -49
rect 161 -51 163 -49
rect 455 -50 457 -48
rect 465 -50 467 -48
rect 759 -50 761 -48
rect 769 -50 771 -48
rect 1064 -50 1066 -48
rect 1074 -50 1076 -48
rect 7 -63 9 -61
rect 17 -63 19 -61
rect 7 -93 9 -67
rect 17 -93 19 -67
rect 151 -81 153 -55
rect 161 -81 163 -55
rect 311 -62 313 -60
rect 321 -62 323 -60
rect 215 -64 217 -62
rect 225 -64 227 -62
rect 151 -87 153 -85
rect 161 -87 163 -85
rect 215 -94 217 -68
rect 225 -94 227 -68
rect 311 -92 313 -66
rect 321 -92 323 -66
rect 455 -80 457 -54
rect 465 -80 467 -54
rect 519 -63 521 -61
rect 529 -63 531 -61
rect 615 -62 617 -60
rect 625 -62 627 -60
rect 455 -86 457 -84
rect 465 -86 467 -84
rect 7 -99 9 -97
rect 17 -99 19 -97
rect 519 -93 521 -67
rect 529 -93 531 -67
rect 615 -92 617 -66
rect 625 -92 627 -66
rect 759 -80 761 -54
rect 769 -80 771 -54
rect 823 -63 825 -61
rect 833 -63 835 -61
rect 920 -62 922 -60
rect 930 -62 932 -60
rect 759 -86 761 -84
rect 769 -86 771 -84
rect 311 -98 313 -96
rect 321 -98 323 -96
rect 823 -93 825 -67
rect 833 -93 835 -67
rect 920 -92 922 -66
rect 930 -92 932 -66
rect 1064 -80 1066 -54
rect 1074 -80 1076 -54
rect 1128 -63 1130 -61
rect 1138 -63 1140 -61
rect 1064 -86 1066 -84
rect 1074 -86 1076 -84
rect 215 -100 217 -98
rect 225 -100 227 -98
rect 519 -99 521 -97
rect 529 -99 531 -97
rect 615 -98 617 -96
rect 625 -98 627 -96
rect 1128 -93 1130 -67
rect 1138 -93 1140 -67
rect 823 -99 825 -97
rect 833 -99 835 -97
rect 920 -98 922 -96
rect 930 -98 932 -96
rect 1128 -99 1130 -97
rect 1138 -99 1140 -97
<< ndiffusion >>
rect -32 -22 -28 -18
rect -26 -22 -22 -18
rect -8 -22 -6 -18
rect -4 -22 6 -18
rect 8 -22 10 -18
rect 22 -22 24 -18
rect 26 -22 32 -18
rect 34 -22 36 -18
rect 48 -22 52 -18
rect 54 -22 58 -18
rect 123 -22 127 -18
rect 129 -22 133 -18
rect 147 -22 149 -18
rect 151 -22 161 -18
rect 163 -22 165 -18
rect 177 -22 179 -18
rect 181 -22 187 -18
rect 189 -22 191 -18
rect 203 -22 207 -18
rect 209 -22 213 -18
rect 272 -21 276 -17
rect 278 -21 282 -17
rect 296 -21 298 -17
rect 300 -21 310 -17
rect 312 -21 314 -17
rect 326 -21 328 -17
rect 330 -21 336 -17
rect 338 -21 340 -17
rect 352 -21 356 -17
rect 358 -21 362 -17
rect 427 -21 431 -17
rect 433 -21 437 -17
rect 451 -21 453 -17
rect 455 -21 465 -17
rect 467 -21 469 -17
rect 481 -21 483 -17
rect 485 -21 491 -17
rect 493 -21 495 -17
rect 507 -21 511 -17
rect 513 -21 517 -17
rect 576 -21 580 -17
rect 582 -21 586 -17
rect 600 -21 602 -17
rect 604 -21 614 -17
rect 616 -21 618 -17
rect 630 -21 632 -17
rect 634 -21 640 -17
rect 642 -21 644 -17
rect 656 -21 660 -17
rect 662 -21 666 -17
rect 731 -21 735 -17
rect 737 -21 741 -17
rect 755 -21 757 -17
rect 759 -21 769 -17
rect 771 -21 773 -17
rect 785 -21 787 -17
rect 789 -21 795 -17
rect 797 -21 799 -17
rect 811 -21 815 -17
rect 817 -21 821 -17
rect 881 -21 885 -17
rect 887 -21 891 -17
rect 905 -21 907 -17
rect 909 -21 919 -17
rect 921 -21 923 -17
rect 935 -21 937 -17
rect 939 -21 945 -17
rect 947 -21 949 -17
rect 961 -21 965 -17
rect 967 -21 971 -17
rect 1036 -21 1040 -17
rect 1042 -21 1046 -17
rect 1060 -21 1062 -17
rect 1064 -21 1074 -17
rect 1076 -21 1078 -17
rect 1090 -21 1092 -17
rect 1094 -21 1100 -17
rect 1102 -21 1104 -17
rect 1116 -21 1120 -17
rect 1122 -21 1126 -17
rect 141 -85 143 -81
rect 147 -85 151 -81
rect 153 -85 161 -81
rect 163 -85 167 -81
rect 171 -85 173 -81
rect -3 -97 -1 -93
rect 3 -97 7 -93
rect 9 -97 17 -93
rect 19 -97 23 -93
rect 27 -97 29 -93
rect 445 -84 447 -80
rect 451 -84 455 -80
rect 457 -84 465 -80
rect 467 -84 471 -80
rect 475 -84 477 -80
rect 205 -98 207 -94
rect 211 -98 215 -94
rect 217 -98 225 -94
rect 227 -98 231 -94
rect 235 -98 237 -94
rect 301 -96 303 -92
rect 307 -96 311 -92
rect 313 -96 321 -92
rect 323 -96 327 -92
rect 331 -96 333 -92
rect 749 -84 751 -80
rect 755 -84 759 -80
rect 761 -84 769 -80
rect 771 -84 775 -80
rect 779 -84 781 -80
rect 509 -97 511 -93
rect 515 -97 519 -93
rect 521 -97 529 -93
rect 531 -97 535 -93
rect 539 -97 541 -93
rect 605 -96 607 -92
rect 611 -96 615 -92
rect 617 -96 625 -92
rect 627 -96 631 -92
rect 635 -96 637 -92
rect 1054 -84 1056 -80
rect 1060 -84 1064 -80
rect 1066 -84 1074 -80
rect 1076 -84 1080 -80
rect 1084 -84 1086 -80
rect 813 -97 815 -93
rect 819 -97 823 -93
rect 825 -97 833 -93
rect 835 -97 839 -93
rect 843 -97 845 -93
rect 910 -96 912 -92
rect 916 -96 920 -92
rect 922 -96 930 -92
rect 932 -96 936 -92
rect 940 -96 942 -92
rect 1118 -97 1120 -93
rect 1124 -97 1128 -93
rect 1130 -97 1138 -93
rect 1140 -97 1144 -93
rect 1148 -97 1150 -93
<< pdiffusion >>
rect -32 10 -28 14
rect -26 10 -22 14
rect -8 10 -6 14
rect -4 10 2 14
rect 4 10 10 14
rect 22 10 24 14
rect 26 10 32 14
rect 34 10 36 14
rect 48 10 52 14
rect 54 10 58 14
rect 123 10 127 14
rect 129 10 133 14
rect 147 10 149 14
rect 151 10 157 14
rect 159 10 165 14
rect 177 10 179 14
rect 181 10 187 14
rect 189 10 191 14
rect 203 10 207 14
rect 209 10 213 14
rect 272 11 276 15
rect 278 11 282 15
rect 296 11 298 15
rect 300 11 306 15
rect 308 11 314 15
rect 326 11 328 15
rect 330 11 336 15
rect 338 11 340 15
rect 352 11 356 15
rect 358 11 362 15
rect 427 11 431 15
rect 433 11 437 15
rect 451 11 453 15
rect 455 11 461 15
rect 463 11 469 15
rect 481 11 483 15
rect 485 11 491 15
rect 493 11 495 15
rect 507 11 511 15
rect 513 11 517 15
rect 576 11 580 15
rect 582 11 586 15
rect 600 11 602 15
rect 604 11 610 15
rect 612 11 618 15
rect 630 11 632 15
rect 634 11 640 15
rect 642 11 644 15
rect 656 11 660 15
rect 662 11 666 15
rect 731 11 735 15
rect 737 11 741 15
rect 755 11 757 15
rect 759 11 765 15
rect 767 11 773 15
rect 785 11 787 15
rect 789 11 795 15
rect 797 11 799 15
rect 811 11 815 15
rect 817 11 821 15
rect 881 11 885 15
rect 887 11 891 15
rect 905 11 907 15
rect 909 11 915 15
rect 917 11 923 15
rect 935 11 937 15
rect 939 11 945 15
rect 947 11 949 15
rect 961 11 965 15
rect 967 11 971 15
rect 1036 11 1040 15
rect 1042 11 1046 15
rect 1060 11 1062 15
rect 1064 11 1070 15
rect 1072 11 1078 15
rect 1090 11 1092 15
rect 1094 11 1100 15
rect 1102 11 1104 15
rect 1116 11 1120 15
rect 1122 11 1126 15
rect 141 -55 143 -51
rect 147 -55 151 -51
rect 153 -55 155 -51
rect 159 -55 161 -51
rect 163 -55 167 -51
rect 171 -55 173 -51
rect 445 -54 447 -50
rect 451 -54 455 -50
rect 457 -54 459 -50
rect 463 -54 465 -50
rect 467 -54 471 -50
rect 475 -54 477 -50
rect 749 -54 751 -50
rect 755 -54 759 -50
rect 761 -54 763 -50
rect 767 -54 769 -50
rect 771 -54 775 -50
rect 779 -54 781 -50
rect 1054 -54 1056 -50
rect 1060 -54 1064 -50
rect 1066 -54 1068 -50
rect 1072 -54 1074 -50
rect 1076 -54 1080 -50
rect 1084 -54 1086 -50
rect -3 -67 -1 -63
rect 3 -67 7 -63
rect 9 -67 11 -63
rect 15 -67 17 -63
rect 19 -67 23 -63
rect 27 -67 29 -63
rect 205 -68 207 -64
rect 211 -68 215 -64
rect 217 -68 219 -64
rect 223 -68 225 -64
rect 227 -68 231 -64
rect 235 -68 237 -64
rect 301 -66 303 -62
rect 307 -66 311 -62
rect 313 -66 315 -62
rect 319 -66 321 -62
rect 323 -66 327 -62
rect 331 -66 333 -62
rect 509 -67 511 -63
rect 515 -67 519 -63
rect 521 -67 523 -63
rect 527 -67 529 -63
rect 531 -67 535 -63
rect 539 -67 541 -63
rect 605 -66 607 -62
rect 611 -66 615 -62
rect 617 -66 619 -62
rect 623 -66 625 -62
rect 627 -66 631 -62
rect 635 -66 637 -62
rect 813 -67 815 -63
rect 819 -67 823 -63
rect 825 -67 827 -63
rect 831 -67 833 -63
rect 835 -67 839 -63
rect 843 -67 845 -63
rect 910 -66 912 -62
rect 916 -66 920 -62
rect 922 -66 924 -62
rect 928 -66 930 -62
rect 932 -66 936 -62
rect 940 -66 942 -62
rect 1118 -67 1120 -63
rect 1124 -67 1128 -63
rect 1130 -67 1132 -63
rect 1136 -67 1138 -63
rect 1140 -67 1144 -63
rect 1148 -67 1150 -63
<< metal1 >>
rect -36 24 -20 28
rect -16 24 14 28
rect 18 24 48 28
rect 52 24 66 28
rect 119 24 135 28
rect 139 24 169 28
rect 173 24 203 28
rect 207 24 221 28
rect 268 25 284 29
rect 288 25 318 29
rect 322 25 352 29
rect 356 25 370 29
rect 423 25 439 29
rect 443 25 473 29
rect 477 25 507 29
rect 511 25 525 29
rect 572 25 588 29
rect 592 25 622 29
rect 626 25 656 29
rect 660 25 674 29
rect 727 25 743 29
rect 747 25 777 29
rect 781 25 811 29
rect 815 25 829 29
rect 877 25 893 29
rect 897 25 927 29
rect 931 25 961 29
rect 965 25 979 29
rect 1032 25 1048 29
rect 1052 25 1082 29
rect 1086 25 1116 29
rect 1120 25 1134 29
rect -36 14 -32 24
rect -12 14 -8 24
rect 36 14 40 24
rect 58 14 62 24
rect -22 6 -18 10
rect -22 2 -10 6
rect -48 -6 -32 -2
rect -48 -73 -44 -6
rect -40 -10 -36 -6
rect -22 -18 -18 2
rect 0 -10 6 -8
rect 0 -12 2 -10
rect 10 -18 14 10
rect 119 14 123 24
rect 143 14 147 24
rect 191 14 195 24
rect 213 14 217 24
rect 18 -18 22 10
rect 44 -8 48 10
rect 133 6 137 10
rect 62 2 110 6
rect 38 -12 48 -8
rect 106 -2 110 2
rect 133 2 145 6
rect 106 -6 123 -2
rect 44 -18 48 -12
rect 58 -14 74 -10
rect -36 -28 -32 -22
rect -12 -28 -8 -22
rect 36 -28 40 -22
rect 58 -28 62 -22
rect -36 -32 -22 -28
rect -18 -32 28 -28
rect 32 -32 46 -28
rect 50 -32 66 -28
rect -5 -59 -1 -55
rect 3 -59 11 -55
rect 15 -59 23 -55
rect 27 -59 31 -55
rect -1 -63 3 -59
rect 23 -63 27 -59
rect 11 -73 15 -67
rect -48 -77 3 -73
rect 11 -77 27 -73
rect -12 -87 13 -83
rect 23 -84 27 -77
rect -12 -108 -8 -87
rect 23 -93 27 -88
rect -1 -101 3 -97
rect -5 -105 -1 -101
rect 3 -105 12 -101
rect 16 -105 23 -101
rect 27 -105 31 -101
rect 70 -108 74 -14
rect 106 -71 110 -6
rect 115 -10 119 -6
rect 133 -18 137 2
rect 155 -10 161 -8
rect 155 -12 157 -10
rect 165 -18 169 10
rect 268 15 272 25
rect 292 15 296 25
rect 340 15 344 25
rect 362 15 366 25
rect 173 -18 177 10
rect 199 -8 203 10
rect 282 7 286 11
rect 218 2 224 6
rect 282 3 294 7
rect 193 -12 203 -8
rect 256 -5 272 -1
rect 199 -18 203 -12
rect 213 -14 230 -10
rect 119 -28 123 -22
rect 143 -28 147 -22
rect 191 -28 195 -22
rect 213 -28 217 -22
rect 119 -32 133 -28
rect 137 -32 183 -28
rect 187 -32 201 -28
rect 205 -32 221 -28
rect 226 -36 230 -14
rect 128 -40 230 -36
rect 128 -61 132 -40
rect 139 -47 143 -43
rect 147 -47 155 -43
rect 159 -47 167 -43
rect 171 -47 175 -43
rect 143 -51 147 -47
rect 167 -51 171 -47
rect 155 -61 159 -55
rect 203 -60 207 -56
rect 211 -60 219 -56
rect 223 -60 231 -56
rect 235 -60 239 -56
rect 128 -65 147 -61
rect 155 -65 171 -61
rect 106 -75 157 -71
rect 167 -74 171 -65
rect 207 -64 211 -60
rect 231 -64 235 -60
rect 219 -74 223 -68
rect 256 -72 260 -5
rect 264 -9 268 -5
rect 282 -17 286 3
rect 304 -9 310 -7
rect 304 -11 306 -9
rect 314 -17 318 11
rect 423 15 427 25
rect 447 15 451 25
rect 495 15 499 25
rect 517 15 521 25
rect 322 -17 326 11
rect 348 -7 352 11
rect 437 7 441 11
rect 366 3 414 7
rect 342 -11 352 -7
rect 410 -1 414 3
rect 437 3 449 7
rect 410 -5 427 -1
rect 348 -17 352 -11
rect 362 -13 378 -9
rect 268 -27 272 -21
rect 292 -27 296 -21
rect 340 -27 344 -21
rect 362 -27 366 -21
rect 268 -31 282 -27
rect 286 -31 332 -27
rect 336 -31 350 -27
rect 354 -31 370 -27
rect 299 -58 303 -54
rect 307 -58 315 -54
rect 319 -58 327 -54
rect 331 -58 335 -54
rect 303 -62 307 -58
rect 327 -62 331 -58
rect 315 -72 319 -66
rect 167 -78 211 -74
rect 219 -78 235 -74
rect 256 -76 307 -72
rect 315 -76 331 -72
rect 167 -81 171 -78
rect 231 -82 235 -78
rect 143 -89 147 -85
rect 204 -88 221 -84
rect 139 -93 143 -89
rect 147 -93 155 -89
rect 159 -93 167 -89
rect 171 -93 175 -89
rect 231 -94 235 -86
rect 292 -86 317 -82
rect 327 -83 331 -76
rect 207 -102 211 -98
rect 203 -106 207 -102
rect 211 -106 219 -102
rect 223 -106 231 -102
rect 235 -106 239 -102
rect -12 -112 74 -108
rect 292 -107 296 -86
rect 327 -92 331 -87
rect 303 -100 307 -96
rect 299 -104 303 -100
rect 307 -104 316 -100
rect 320 -104 327 -100
rect 331 -104 335 -100
rect 374 -107 378 -13
rect 410 -70 414 -5
rect 419 -9 423 -5
rect 437 -17 441 3
rect 459 -9 465 -7
rect 459 -11 461 -9
rect 469 -17 473 11
rect 572 15 576 25
rect 596 15 600 25
rect 644 15 648 25
rect 666 15 670 25
rect 477 -17 481 11
rect 503 -7 507 11
rect 586 7 590 11
rect 522 3 528 7
rect 586 3 598 7
rect 497 -11 507 -7
rect 560 -5 576 -1
rect 503 -17 507 -11
rect 517 -13 534 -9
rect 423 -27 427 -21
rect 447 -27 451 -21
rect 495 -27 499 -21
rect 517 -27 521 -21
rect 423 -31 437 -27
rect 441 -31 487 -27
rect 491 -31 505 -27
rect 509 -31 525 -27
rect 530 -35 534 -13
rect 432 -39 534 -35
rect 432 -40 436 -39
rect 432 -60 436 -44
rect 443 -46 447 -42
rect 451 -46 459 -42
rect 463 -46 471 -42
rect 475 -46 479 -42
rect 447 -50 451 -46
rect 471 -50 475 -46
rect 459 -60 463 -54
rect 507 -59 511 -55
rect 515 -59 523 -55
rect 527 -59 535 -55
rect 539 -59 543 -55
rect 432 -64 451 -60
rect 459 -64 475 -60
rect 410 -74 461 -70
rect 471 -73 475 -64
rect 511 -63 515 -59
rect 535 -63 539 -59
rect 523 -73 527 -67
rect 560 -72 564 -5
rect 568 -9 572 -5
rect 586 -17 590 3
rect 608 -9 614 -7
rect 608 -11 610 -9
rect 618 -17 622 11
rect 727 15 731 25
rect 751 15 755 25
rect 799 15 803 25
rect 821 15 825 25
rect 626 -17 630 11
rect 652 -7 656 11
rect 741 7 745 11
rect 670 3 718 7
rect 646 -11 656 -7
rect 714 -1 718 3
rect 741 3 753 7
rect 714 -5 731 -1
rect 652 -17 656 -11
rect 666 -13 682 -9
rect 572 -27 576 -21
rect 596 -27 600 -21
rect 644 -27 648 -21
rect 666 -27 670 -21
rect 572 -31 586 -27
rect 590 -31 636 -27
rect 640 -31 654 -27
rect 658 -31 674 -27
rect 603 -58 607 -54
rect 611 -58 619 -54
rect 623 -58 631 -54
rect 635 -58 639 -54
rect 607 -62 611 -58
rect 631 -62 635 -58
rect 619 -72 623 -66
rect 471 -77 515 -73
rect 523 -77 539 -73
rect 560 -76 611 -72
rect 619 -76 635 -72
rect 471 -80 475 -77
rect 535 -80 539 -77
rect 447 -88 451 -84
rect 508 -87 525 -83
rect 443 -92 447 -88
rect 451 -92 459 -88
rect 463 -92 471 -88
rect 475 -92 479 -88
rect 535 -93 539 -84
rect 596 -86 621 -82
rect 631 -83 635 -76
rect 511 -101 515 -97
rect 507 -105 511 -101
rect 515 -105 523 -101
rect 527 -105 535 -101
rect 539 -105 543 -101
rect 292 -111 378 -107
rect 596 -107 600 -86
rect 631 -92 635 -87
rect 607 -100 611 -96
rect 603 -104 607 -100
rect 611 -104 620 -100
rect 624 -104 631 -100
rect 635 -104 639 -100
rect 678 -107 682 -13
rect 714 -70 718 -5
rect 723 -9 727 -5
rect 741 -17 745 3
rect 763 -9 769 -7
rect 763 -11 765 -9
rect 773 -17 777 11
rect 877 15 881 25
rect 901 15 905 25
rect 949 15 953 25
rect 971 15 975 25
rect 781 -17 785 11
rect 807 -7 811 11
rect 891 7 895 11
rect 826 3 832 7
rect 891 3 903 7
rect 801 -11 811 -7
rect 865 -5 881 -1
rect 807 -17 811 -11
rect 821 -13 838 -9
rect 727 -27 731 -21
rect 751 -27 755 -21
rect 799 -27 803 -21
rect 821 -27 825 -21
rect 727 -31 741 -27
rect 745 -31 791 -27
rect 795 -31 809 -27
rect 813 -31 829 -27
rect 834 -35 838 -13
rect 736 -36 838 -35
rect 740 -39 838 -36
rect 736 -60 740 -40
rect 747 -46 751 -42
rect 755 -46 763 -42
rect 767 -46 775 -42
rect 779 -46 783 -42
rect 751 -50 755 -46
rect 775 -50 779 -46
rect 763 -60 767 -54
rect 811 -59 815 -55
rect 819 -59 827 -55
rect 831 -59 839 -55
rect 843 -59 847 -55
rect 736 -64 755 -60
rect 763 -64 779 -60
rect 714 -74 765 -70
rect 775 -73 779 -64
rect 815 -63 819 -59
rect 839 -63 843 -59
rect 827 -73 831 -67
rect 865 -72 869 -5
rect 873 -9 877 -5
rect 891 -17 895 3
rect 913 -9 919 -7
rect 913 -11 915 -9
rect 923 -17 927 11
rect 1032 15 1036 25
rect 1056 15 1060 25
rect 1104 15 1108 25
rect 1126 15 1130 25
rect 931 -17 935 11
rect 957 -7 961 11
rect 1046 7 1050 11
rect 975 3 1023 7
rect 951 -11 961 -7
rect 1019 -1 1023 3
rect 1046 3 1058 7
rect 1019 -5 1036 -1
rect 957 -17 961 -11
rect 971 -13 987 -9
rect 877 -27 881 -21
rect 901 -27 905 -21
rect 949 -27 953 -21
rect 971 -27 975 -21
rect 877 -31 891 -27
rect 895 -31 941 -27
rect 945 -31 959 -27
rect 963 -31 979 -27
rect 908 -58 912 -54
rect 916 -58 924 -54
rect 928 -58 936 -54
rect 940 -58 944 -54
rect 912 -62 916 -58
rect 936 -62 940 -58
rect 924 -72 928 -66
rect 775 -77 819 -73
rect 827 -77 843 -73
rect 865 -76 916 -72
rect 924 -76 940 -72
rect 775 -80 779 -77
rect 839 -82 843 -77
rect 751 -88 755 -84
rect 812 -87 829 -83
rect 747 -92 751 -88
rect 755 -92 763 -88
rect 767 -92 775 -88
rect 779 -92 783 -88
rect 839 -93 843 -86
rect 901 -86 926 -82
rect 936 -83 940 -76
rect 815 -101 819 -97
rect 811 -105 815 -101
rect 819 -105 827 -101
rect 831 -105 839 -101
rect 843 -105 847 -101
rect 596 -111 682 -107
rect 901 -107 905 -86
rect 936 -92 940 -87
rect 912 -100 916 -96
rect 908 -104 912 -100
rect 916 -104 925 -100
rect 929 -104 936 -100
rect 940 -104 944 -100
rect 983 -107 987 -13
rect 1019 -70 1023 -5
rect 1028 -9 1032 -5
rect 1046 -17 1050 3
rect 1068 -9 1074 -7
rect 1068 -11 1070 -9
rect 1078 -17 1082 11
rect 1086 -17 1090 11
rect 1112 -7 1116 11
rect 1131 3 1137 7
rect 1106 -11 1116 -7
rect 1112 -17 1116 -11
rect 1126 -13 1143 -9
rect 1032 -27 1036 -21
rect 1056 -27 1060 -21
rect 1104 -27 1108 -21
rect 1126 -27 1130 -21
rect 1032 -31 1046 -27
rect 1050 -31 1096 -27
rect 1100 -31 1114 -27
rect 1118 -31 1134 -27
rect 1139 -35 1143 -13
rect 1041 -38 1143 -35
rect 1045 -39 1143 -38
rect 1041 -60 1045 -42
rect 1052 -46 1056 -42
rect 1060 -46 1068 -42
rect 1072 -46 1080 -42
rect 1084 -46 1088 -42
rect 1056 -50 1060 -46
rect 1080 -50 1084 -46
rect 1068 -60 1072 -54
rect 1116 -59 1120 -55
rect 1124 -59 1132 -55
rect 1136 -59 1144 -55
rect 1148 -59 1152 -55
rect 1041 -64 1060 -60
rect 1068 -64 1084 -60
rect 1019 -74 1070 -70
rect 1080 -73 1084 -64
rect 1120 -63 1124 -59
rect 1144 -63 1148 -59
rect 1132 -73 1136 -67
rect 1080 -77 1124 -73
rect 1132 -77 1148 -73
rect 1080 -80 1084 -77
rect 1056 -88 1060 -84
rect 1117 -87 1134 -83
rect 1052 -92 1056 -88
rect 1060 -92 1068 -88
rect 1072 -92 1080 -88
rect 1084 -92 1088 -88
rect 1144 -93 1148 -77
rect 1120 -101 1124 -97
rect 1116 -105 1120 -101
rect 1124 -105 1132 -101
rect 1136 -105 1144 -101
rect 1148 -105 1152 -101
rect 901 -111 987 -107
<< metal2 >>
rect 18 2 58 6
rect 173 2 214 6
rect 322 3 362 7
rect 477 3 518 7
rect 626 3 666 7
rect 781 3 822 7
rect 931 3 971 7
rect 1086 3 1127 7
rect -12 -10 -4 -8
rect -36 -12 -4 -10
rect 143 -10 151 -8
rect -36 -14 -8 -12
rect 119 -12 151 -10
rect 292 -9 300 -7
rect 119 -14 147 -12
rect 268 -11 300 -9
rect 447 -9 455 -7
rect 268 -13 296 -11
rect 423 -11 455 -9
rect 596 -9 604 -7
rect 423 -13 451 -11
rect 572 -11 604 -9
rect 751 -9 759 -7
rect 572 -13 600 -11
rect 727 -11 759 -9
rect 901 -9 909 -7
rect 727 -13 755 -11
rect 877 -11 909 -9
rect 1056 -9 1064 -7
rect 877 -13 905 -11
rect 1032 -11 1064 -9
rect 1032 -13 1060 -11
rect 550 -40 736 -36
rect 246 -44 432 -40
rect 246 -82 250 -44
rect 550 -80 554 -40
rect 27 -88 110 -84
rect 106 -98 110 -88
rect 192 -88 200 -84
rect 235 -86 250 -82
rect 331 -87 414 -83
rect 192 -98 196 -88
rect 106 -102 196 -98
rect 410 -97 414 -87
rect 496 -87 504 -83
rect 539 -84 554 -80
rect 856 -42 1041 -38
rect 856 -82 860 -42
rect 635 -87 718 -83
rect 496 -97 500 -87
rect 410 -101 500 -97
rect 714 -97 718 -87
rect 800 -87 808 -83
rect 843 -86 860 -82
rect 940 -87 1023 -83
rect 800 -97 804 -87
rect 714 -101 804 -97
rect 1019 -97 1023 -87
rect 1105 -87 1113 -83
rect 1105 -97 1109 -87
rect 1019 -101 1109 -97
<< ntransistor >>
rect -28 -22 -26 -18
rect -6 -22 -4 -18
rect 6 -22 8 -18
rect 24 -22 26 -18
rect 32 -22 34 -18
rect 52 -22 54 -18
rect 127 -22 129 -18
rect 149 -22 151 -18
rect 161 -22 163 -18
rect 179 -22 181 -18
rect 187 -22 189 -18
rect 207 -22 209 -18
rect 276 -21 278 -17
rect 298 -21 300 -17
rect 310 -21 312 -17
rect 328 -21 330 -17
rect 336 -21 338 -17
rect 356 -21 358 -17
rect 431 -21 433 -17
rect 453 -21 455 -17
rect 465 -21 467 -17
rect 483 -21 485 -17
rect 491 -21 493 -17
rect 511 -21 513 -17
rect 580 -21 582 -17
rect 602 -21 604 -17
rect 614 -21 616 -17
rect 632 -21 634 -17
rect 640 -21 642 -17
rect 660 -21 662 -17
rect 735 -21 737 -17
rect 757 -21 759 -17
rect 769 -21 771 -17
rect 787 -21 789 -17
rect 795 -21 797 -17
rect 815 -21 817 -17
rect 885 -21 887 -17
rect 907 -21 909 -17
rect 919 -21 921 -17
rect 937 -21 939 -17
rect 945 -21 947 -17
rect 965 -21 967 -17
rect 1040 -21 1042 -17
rect 1062 -21 1064 -17
rect 1074 -21 1076 -17
rect 1092 -21 1094 -17
rect 1100 -21 1102 -17
rect 1120 -21 1122 -17
rect 151 -85 153 -81
rect 161 -85 163 -81
rect 7 -97 9 -93
rect 17 -97 19 -93
rect 455 -84 457 -80
rect 465 -84 467 -80
rect 215 -98 217 -94
rect 225 -98 227 -94
rect 311 -96 313 -92
rect 321 -96 323 -92
rect 759 -84 761 -80
rect 769 -84 771 -80
rect 519 -97 521 -93
rect 529 -97 531 -93
rect 615 -96 617 -92
rect 625 -96 627 -92
rect 1064 -84 1066 -80
rect 1074 -84 1076 -80
rect 823 -97 825 -93
rect 833 -97 835 -93
rect 920 -96 922 -92
rect 930 -96 932 -92
rect 1128 -97 1130 -93
rect 1138 -97 1140 -93
<< ptransistor >>
rect -28 10 -26 14
rect -6 10 -4 14
rect 2 10 4 14
rect 24 10 26 14
rect 32 10 34 14
rect 52 10 54 14
rect 127 10 129 14
rect 149 10 151 14
rect 157 10 159 14
rect 179 10 181 14
rect 187 10 189 14
rect 207 10 209 14
rect 276 11 278 15
rect 298 11 300 15
rect 306 11 308 15
rect 328 11 330 15
rect 336 11 338 15
rect 356 11 358 15
rect 431 11 433 15
rect 453 11 455 15
rect 461 11 463 15
rect 483 11 485 15
rect 491 11 493 15
rect 511 11 513 15
rect 580 11 582 15
rect 602 11 604 15
rect 610 11 612 15
rect 632 11 634 15
rect 640 11 642 15
rect 660 11 662 15
rect 735 11 737 15
rect 757 11 759 15
rect 765 11 767 15
rect 787 11 789 15
rect 795 11 797 15
rect 815 11 817 15
rect 885 11 887 15
rect 907 11 909 15
rect 915 11 917 15
rect 937 11 939 15
rect 945 11 947 15
rect 965 11 967 15
rect 1040 11 1042 15
rect 1062 11 1064 15
rect 1070 11 1072 15
rect 1092 11 1094 15
rect 1100 11 1102 15
rect 1120 11 1122 15
rect 151 -55 153 -51
rect 161 -55 163 -51
rect 455 -54 457 -50
rect 465 -54 467 -50
rect 759 -54 761 -50
rect 769 -54 771 -50
rect 1064 -54 1066 -50
rect 1074 -54 1076 -50
rect 7 -67 9 -63
rect 17 -67 19 -63
rect 215 -68 217 -64
rect 225 -68 227 -64
rect 311 -66 313 -62
rect 321 -66 323 -62
rect 519 -67 521 -63
rect 529 -67 531 -63
rect 615 -66 617 -62
rect 625 -66 627 -62
rect 823 -67 825 -63
rect 833 -67 835 -63
rect 920 -66 922 -62
rect 930 -66 932 -62
rect 1128 -67 1130 -63
rect 1138 -67 1140 -63
<< polycontact >>
rect -32 -6 -28 -2
rect -10 2 -6 6
rect 2 -14 6 -10
rect 34 -12 38 -8
rect 123 -6 127 -2
rect 54 -14 58 -10
rect 145 2 149 6
rect 157 -14 161 -10
rect 189 -12 193 -8
rect 272 -5 276 -1
rect 209 -14 213 -10
rect 294 3 298 7
rect 306 -13 310 -9
rect 338 -11 342 -7
rect 427 -5 431 -1
rect 358 -13 362 -9
rect 449 3 453 7
rect 461 -13 465 -9
rect 493 -11 497 -7
rect 576 -5 580 -1
rect 513 -13 517 -9
rect 598 3 602 7
rect 610 -13 614 -9
rect 642 -11 646 -7
rect 731 -5 735 -1
rect 662 -13 666 -9
rect 753 3 757 7
rect 765 -13 769 -9
rect 797 -11 801 -7
rect 881 -5 885 -1
rect 817 -13 821 -9
rect 903 3 907 7
rect 915 -13 919 -9
rect 947 -11 951 -7
rect 1036 -5 1040 -1
rect 967 -13 971 -9
rect 1058 3 1062 7
rect 1070 -13 1074 -9
rect 1102 -11 1106 -7
rect 1122 -13 1126 -9
rect 147 -65 151 -61
rect 3 -77 7 -73
rect 13 -87 17 -83
rect 157 -75 161 -71
rect 451 -64 455 -60
rect 211 -78 215 -74
rect 221 -88 225 -84
rect 307 -76 311 -72
rect 317 -86 321 -82
rect 461 -74 465 -70
rect 755 -64 759 -60
rect 515 -77 519 -73
rect 525 -87 529 -83
rect 611 -76 615 -72
rect 621 -86 625 -82
rect 765 -74 769 -70
rect 1060 -64 1064 -60
rect 819 -77 823 -73
rect 829 -87 833 -83
rect 916 -76 920 -72
rect 926 -86 930 -82
rect 1070 -74 1074 -70
rect 1124 -77 1128 -73
rect 1134 -87 1138 -83
<< ndcontact >>
rect -36 -22 -32 -18
rect -22 -22 -18 -18
rect -12 -22 -8 -18
rect 10 -22 14 -18
rect 18 -22 22 -18
rect 36 -22 40 -18
rect 44 -22 48 -18
rect 58 -22 62 -18
rect 119 -22 123 -18
rect 133 -22 137 -18
rect 143 -22 147 -18
rect 165 -22 169 -18
rect 173 -22 177 -18
rect 191 -22 195 -18
rect 199 -22 203 -18
rect 213 -22 217 -18
rect 268 -21 272 -17
rect 282 -21 286 -17
rect 292 -21 296 -17
rect 314 -21 318 -17
rect 322 -21 326 -17
rect 340 -21 344 -17
rect 348 -21 352 -17
rect 362 -21 366 -17
rect 423 -21 427 -17
rect 437 -21 441 -17
rect 447 -21 451 -17
rect 469 -21 473 -17
rect 477 -21 481 -17
rect 495 -21 499 -17
rect 503 -21 507 -17
rect 517 -21 521 -17
rect 572 -21 576 -17
rect 586 -21 590 -17
rect 596 -21 600 -17
rect 618 -21 622 -17
rect 626 -21 630 -17
rect 644 -21 648 -17
rect 652 -21 656 -17
rect 666 -21 670 -17
rect 727 -21 731 -17
rect 741 -21 745 -17
rect 751 -21 755 -17
rect 773 -21 777 -17
rect 781 -21 785 -17
rect 799 -21 803 -17
rect 807 -21 811 -17
rect 821 -21 825 -17
rect 877 -21 881 -17
rect 891 -21 895 -17
rect 901 -21 905 -17
rect 923 -21 927 -17
rect 931 -21 935 -17
rect 949 -21 953 -17
rect 957 -21 961 -17
rect 971 -21 975 -17
rect 1032 -21 1036 -17
rect 1046 -21 1050 -17
rect 1056 -21 1060 -17
rect 1078 -21 1082 -17
rect 1086 -21 1090 -17
rect 1104 -21 1108 -17
rect 1112 -21 1116 -17
rect 1126 -21 1130 -17
rect 143 -85 147 -81
rect 167 -85 171 -81
rect -1 -97 3 -93
rect 23 -97 27 -93
rect 447 -84 451 -80
rect 471 -84 475 -80
rect 207 -98 211 -94
rect 231 -98 235 -94
rect 303 -96 307 -92
rect 327 -96 331 -92
rect 751 -84 755 -80
rect 775 -84 779 -80
rect 511 -97 515 -93
rect 535 -97 539 -93
rect 607 -96 611 -92
rect 631 -96 635 -92
rect 1056 -84 1060 -80
rect 1080 -84 1084 -80
rect 815 -97 819 -93
rect 839 -97 843 -93
rect 912 -96 916 -92
rect 936 -96 940 -92
rect 1120 -97 1124 -93
rect 1144 -97 1148 -93
<< pdcontact >>
rect -36 10 -32 14
rect -22 10 -18 14
rect -12 10 -8 14
rect 10 10 14 14
rect 18 10 22 14
rect 36 10 40 14
rect 44 10 48 14
rect 58 10 62 14
rect 119 10 123 14
rect 133 10 137 14
rect 143 10 147 14
rect 165 10 169 14
rect 173 10 177 14
rect 191 10 195 14
rect 199 10 203 14
rect 213 10 217 14
rect 268 11 272 15
rect 282 11 286 15
rect 292 11 296 15
rect 314 11 318 15
rect 322 11 326 15
rect 340 11 344 15
rect 348 11 352 15
rect 362 11 366 15
rect 423 11 427 15
rect 437 11 441 15
rect 447 11 451 15
rect 469 11 473 15
rect 477 11 481 15
rect 495 11 499 15
rect 503 11 507 15
rect 517 11 521 15
rect 572 11 576 15
rect 586 11 590 15
rect 596 11 600 15
rect 618 11 622 15
rect 626 11 630 15
rect 644 11 648 15
rect 652 11 656 15
rect 666 11 670 15
rect 727 11 731 15
rect 741 11 745 15
rect 751 11 755 15
rect 773 11 777 15
rect 781 11 785 15
rect 799 11 803 15
rect 807 11 811 15
rect 821 11 825 15
rect 877 11 881 15
rect 891 11 895 15
rect 901 11 905 15
rect 923 11 927 15
rect 931 11 935 15
rect 949 11 953 15
rect 957 11 961 15
rect 971 11 975 15
rect 1032 11 1036 15
rect 1046 11 1050 15
rect 1056 11 1060 15
rect 1078 11 1082 15
rect 1086 11 1090 15
rect 1104 11 1108 15
rect 1112 11 1116 15
rect 1126 11 1130 15
rect 143 -55 147 -51
rect 155 -55 159 -51
rect 167 -55 171 -51
rect 447 -54 451 -50
rect 459 -54 463 -50
rect 471 -54 475 -50
rect 751 -54 755 -50
rect 763 -54 767 -50
rect 775 -54 779 -50
rect 1056 -54 1060 -50
rect 1068 -54 1072 -50
rect 1080 -54 1084 -50
rect -1 -67 3 -63
rect 11 -67 15 -63
rect 23 -67 27 -63
rect 207 -68 211 -64
rect 219 -68 223 -64
rect 231 -68 235 -64
rect 303 -66 307 -62
rect 315 -66 319 -62
rect 327 -66 331 -62
rect 511 -67 515 -63
rect 523 -67 527 -63
rect 535 -67 539 -63
rect 607 -66 611 -62
rect 619 -66 623 -62
rect 631 -66 635 -62
rect 815 -67 819 -63
rect 827 -67 831 -63
rect 839 -67 843 -63
rect 912 -66 916 -62
rect 924 -66 928 -62
rect 936 -66 940 -62
rect 1120 -67 1124 -63
rect 1132 -67 1136 -63
rect 1144 -67 1148 -63
<< m2contact >>
rect -40 -14 -36 -10
rect -4 -12 0 -8
rect 14 2 18 6
rect 58 2 62 6
rect 23 -88 27 -84
rect 115 -14 119 -10
rect 151 -12 155 -8
rect 169 2 173 6
rect 214 2 218 6
rect 264 -13 268 -9
rect 300 -11 304 -7
rect 318 3 322 7
rect 362 3 366 7
rect 200 -88 204 -84
rect 231 -86 235 -82
rect 327 -87 331 -83
rect 419 -13 423 -9
rect 455 -11 459 -7
rect 473 3 477 7
rect 518 3 522 7
rect 432 -44 436 -40
rect 568 -13 572 -9
rect 604 -11 608 -7
rect 622 3 626 7
rect 666 3 670 7
rect 504 -87 508 -83
rect 535 -84 539 -80
rect 631 -87 635 -83
rect 723 -13 727 -9
rect 759 -11 763 -7
rect 777 3 781 7
rect 822 3 826 7
rect 736 -40 740 -36
rect 873 -13 877 -9
rect 909 -11 913 -7
rect 927 3 931 7
rect 971 3 975 7
rect 808 -87 812 -83
rect 839 -86 843 -82
rect 936 -87 940 -83
rect 1028 -13 1032 -9
rect 1064 -11 1068 -7
rect 1082 3 1086 7
rect 1127 3 1131 7
rect 1041 -42 1045 -38
rect 1113 -87 1117 -83
<< psubstratepcontact >>
rect -22 -32 -18 -28
rect 28 -32 32 -28
rect 46 -32 50 -28
rect 133 -32 137 -28
rect 183 -32 187 -28
rect 201 -32 205 -28
rect 282 -31 286 -27
rect 332 -31 336 -27
rect 350 -31 354 -27
rect 437 -31 441 -27
rect 487 -31 491 -27
rect 505 -31 509 -27
rect 586 -31 590 -27
rect 636 -31 640 -27
rect 654 -31 658 -27
rect 741 -31 745 -27
rect 791 -31 795 -27
rect 809 -31 813 -27
rect 891 -31 895 -27
rect 941 -31 945 -27
rect 959 -31 963 -27
rect 1046 -31 1050 -27
rect 1096 -31 1100 -27
rect 1114 -31 1118 -27
rect 143 -93 147 -89
rect 155 -93 159 -89
rect 167 -93 171 -89
rect 447 -92 451 -88
rect 459 -92 463 -88
rect 471 -92 475 -88
rect 751 -92 755 -88
rect 763 -92 767 -88
rect 775 -92 779 -88
rect 1056 -92 1060 -88
rect 1068 -92 1072 -88
rect 1080 -92 1084 -88
rect -1 -105 3 -101
rect 12 -105 16 -101
rect 23 -105 27 -101
rect 207 -106 211 -102
rect 219 -106 223 -102
rect 231 -106 235 -102
rect 303 -104 307 -100
rect 316 -104 320 -100
rect 327 -104 331 -100
rect 511 -105 515 -101
rect 523 -105 527 -101
rect 535 -105 539 -101
rect 607 -104 611 -100
rect 620 -104 624 -100
rect 631 -104 635 -100
rect 815 -105 819 -101
rect 827 -105 831 -101
rect 839 -105 843 -101
rect 912 -104 916 -100
rect 925 -104 929 -100
rect 936 -104 940 -100
rect 1120 -105 1124 -101
rect 1132 -105 1136 -101
rect 1144 -105 1148 -101
<< nsubstratencontact >>
rect -20 24 -16 28
rect 14 24 18 28
rect 48 24 52 28
rect 135 24 139 28
rect 169 24 173 28
rect 203 24 207 28
rect 284 25 288 29
rect 318 25 322 29
rect 352 25 356 29
rect 439 25 443 29
rect 473 25 477 29
rect 507 25 511 29
rect 588 25 592 29
rect 622 25 626 29
rect 656 25 660 29
rect 743 25 747 29
rect 777 25 781 29
rect 811 25 815 29
rect 893 25 897 29
rect 927 25 931 29
rect 961 25 965 29
rect 1048 25 1052 29
rect 1082 25 1086 29
rect 1116 25 1120 29
rect 143 -47 147 -43
rect 155 -47 159 -43
rect 167 -47 171 -43
rect 447 -46 451 -42
rect 459 -46 463 -42
rect 471 -46 475 -42
rect 751 -46 755 -42
rect 763 -46 767 -42
rect 775 -46 779 -42
rect 1056 -46 1060 -42
rect 1068 -46 1072 -42
rect 1080 -46 1084 -42
rect -1 -59 3 -55
rect 11 -59 15 -55
rect 23 -59 27 -55
rect 207 -60 211 -56
rect 219 -60 223 -56
rect 231 -60 235 -56
rect 303 -58 307 -54
rect 315 -58 319 -54
rect 327 -58 331 -54
rect 511 -59 515 -55
rect 523 -59 527 -55
rect 535 -59 539 -55
rect 607 -58 611 -54
rect 619 -58 623 -54
rect 631 -58 635 -54
rect 815 -59 819 -55
rect 827 -59 831 -55
rect 839 -59 843 -55
rect 912 -58 916 -54
rect 924 -58 928 -54
rect 936 -58 940 -54
rect 1120 -59 1124 -55
rect 1132 -59 1136 -55
rect 1144 -59 1148 -55
<< labels >>
rlabel metal1 4 25 6 27 5 VDD
rlabel metal1 8 -31 10 -29 1 GND
rlabel metal1 159 25 161 27 5 VDD
rlabel metal1 163 -31 165 -29 1 GND
rlabel nsubstratencontact 156 -46 158 -44 1 VDD
rlabel psubstratepcontact 156 -92 158 -90 1 GND
rlabel nsubstratencontact 12 -58 14 -56 1 VDD
rlabel psubstratepcontact 12 -104 14 -102 1 GND
rlabel nsubstratencontact 220 -59 222 -57 1 VDD
rlabel psubstratepcontact 220 -105 222 -103 1 GND
rlabel metal1 129 -39 131 -37 1 Cin
rlabel metal1 308 26 310 28 5 VDD
rlabel metal1 312 -30 314 -28 1 GND
rlabel metal1 463 26 465 28 5 VDD
rlabel metal1 467 -30 469 -28 1 GND
rlabel nsubstratencontact 460 -45 462 -43 1 VDD
rlabel psubstratepcontact 460 -91 462 -89 1 GND
rlabel nsubstratencontact 316 -57 318 -55 1 VDD
rlabel psubstratepcontact 316 -103 318 -101 1 GND
rlabel nsubstratencontact 524 -58 526 -56 1 VDD
rlabel psubstratepcontact 524 -104 526 -102 1 GND
rlabel metal1 612 26 614 28 5 VDD
rlabel metal1 616 -30 618 -28 1 GND
rlabel metal1 767 26 769 28 5 VDD
rlabel metal1 771 -30 773 -28 1 GND
rlabel nsubstratencontact 764 -45 766 -43 1 VDD
rlabel psubstratepcontact 764 -91 766 -89 1 GND
rlabel nsubstratencontact 620 -57 622 -55 1 VDD
rlabel psubstratepcontact 620 -103 622 -101 1 GND
rlabel nsubstratencontact 828 -58 830 -56 1 VDD
rlabel psubstratepcontact 828 -104 830 -102 1 GND
rlabel metal1 917 26 919 28 5 VDD
rlabel metal1 921 -30 923 -28 1 GND
rlabel metal1 1072 26 1074 28 5 VDD
rlabel metal1 1076 -30 1078 -28 1 GND
rlabel nsubstratencontact 1069 -45 1071 -43 1 VDD
rlabel psubstratepcontact 1069 -91 1071 -89 1 GND
rlabel nsubstratencontact 925 -57 927 -55 1 VDD
rlabel psubstratepcontact 925 -103 927 -101 1 GND
rlabel nsubstratencontact 1133 -58 1135 -56 1 VDD
rlabel psubstratepcontact 1133 -104 1135 -102 1 GND
rlabel metal1 1145 -76 1147 -74 1 Cout
rlabel polycontact -31 -5 -29 -3 1 A0
rlabel polycontact 55 -13 57 -11 1 B0
rlabel metal1 221 3 223 5 1 S0
rlabel polycontact 273 -4 275 -2 1 A1
rlabel polycontact 359 -12 361 -10 1 B1
rlabel metal1 525 4 527 6 1 S1
rlabel polycontact 577 -4 579 -2 1 A2
rlabel polycontact 663 -12 665 -10 1 B2
rlabel metal1 829 4 831 6 1 S2
rlabel polycontact 882 -4 884 -2 1 A3
rlabel polycontact 968 -12 970 -10 1 B3
rlabel metal1 1134 4 1136 6 1 S3
<< end >>
