magic
tech scmos
timestamp 1461798863
<< nwell >>
rect -40 8 70 30
<< polysilicon >>
rect 2 20 54 22
rect -28 14 -26 16
rect -6 14 -4 16
rect 2 14 4 20
rect 24 14 26 16
rect 32 14 34 16
rect 52 14 54 20
rect -28 -18 -26 10
rect -6 2 -4 10
rect -16 0 -4 2
rect -28 -24 -26 -22
rect -16 -26 -14 0
rect 2 -2 4 10
rect -8 -4 4 -2
rect -8 -14 -6 -4
rect 24 -10 26 10
rect 6 -12 26 -10
rect -8 -16 -4 -14
rect -6 -18 -4 -16
rect 6 -18 8 -12
rect 24 -18 26 -16
rect 32 -18 34 10
rect 52 -18 54 10
rect -6 -24 -4 -22
rect 6 -24 8 -22
rect 24 -26 26 -22
rect 32 -24 34 -22
rect 52 -24 54 -22
rect -16 -28 26 -26
<< ndiffusion >>
rect -32 -22 -28 -18
rect -26 -22 -22 -18
rect -8 -22 -6 -18
rect -4 -22 6 -18
rect 8 -22 10 -18
rect 22 -22 24 -18
rect 26 -22 32 -18
rect 34 -22 36 -18
rect 48 -22 52 -18
rect 54 -22 58 -18
<< pdiffusion >>
rect -32 10 -28 14
rect -26 10 -22 14
rect -8 10 -6 14
rect -4 10 2 14
rect 4 10 10 14
rect 22 10 24 14
rect 26 10 32 14
rect 34 10 36 14
rect 48 10 52 14
rect 54 10 58 14
<< metal1 >>
rect -36 24 -20 28
rect -16 24 14 28
rect 18 24 48 28
rect 52 24 66 28
rect -36 14 -32 24
rect -12 14 -8 24
rect 36 14 40 24
rect 58 14 62 24
rect -22 6 -18 10
rect -22 2 -10 6
rect -40 -6 -32 -2
rect -40 -10 -36 -6
rect -22 -18 -18 2
rect 0 -10 6 -8
rect 0 -12 2 -10
rect 10 -18 14 10
rect 18 -18 22 10
rect 44 -8 48 10
rect 62 2 66 6
rect 38 -12 48 -8
rect 44 -18 48 -12
rect 58 -14 66 -10
rect -36 -28 -32 -22
rect -12 -28 -8 -22
rect 36 -28 40 -22
rect 58 -28 62 -22
rect -36 -32 -22 -28
rect -18 -32 28 -28
rect 32 -32 46 -28
rect 50 -32 66 -28
<< metal2 >>
rect 18 2 58 6
rect -12 -10 -4 -8
rect -36 -12 -4 -10
rect -36 -14 -8 -12
<< ntransistor >>
rect -28 -22 -26 -18
rect -6 -22 -4 -18
rect 6 -22 8 -18
rect 24 -22 26 -18
rect 32 -22 34 -18
rect 52 -22 54 -18
<< ptransistor >>
rect -28 10 -26 14
rect -6 10 -4 14
rect 2 10 4 14
rect 24 10 26 14
rect 32 10 34 14
rect 52 10 54 14
<< polycontact >>
rect -32 -6 -28 -2
rect -10 2 -6 6
rect 2 -14 6 -10
rect 34 -12 38 -8
rect 54 -14 58 -10
<< ndcontact >>
rect -36 -22 -32 -18
rect -22 -22 -18 -18
rect -12 -22 -8 -18
rect 10 -22 14 -18
rect 18 -22 22 -18
rect 36 -22 40 -18
rect 44 -22 48 -18
rect 58 -22 62 -18
<< pdcontact >>
rect -36 10 -32 14
rect -22 10 -18 14
rect -12 10 -8 14
rect 10 10 14 14
rect 18 10 22 14
rect 36 10 40 14
rect 44 10 48 14
rect 58 10 62 14
<< m2contact >>
rect -40 -14 -36 -10
rect -4 -12 0 -8
rect 14 2 18 6
rect 58 2 62 6
<< psubstratepcontact >>
rect -22 -32 -18 -28
rect 28 -32 32 -28
rect 46 -32 50 -28
<< nsubstratencontact >>
rect -20 24 -16 28
rect 14 24 18 28
rect 48 24 52 28
<< labels >>
rlabel polycontact -30 -5 -28 -3 1 A
rlabel polycontact 54 -13 56 -11 1 B
rlabel m2contact 59 3 61 5 1 Y
rlabel metal1 4 25 6 27 5 VDD
rlabel metal1 8 -31 10 -29 1 GND
<< end >>
